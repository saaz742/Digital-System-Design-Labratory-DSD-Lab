`timescale 1ns / 1ps

module testdiv;

	// Instantiate the Unit Under Test (UUT)
	div uut (
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

